----------------------------------------------------------------------------------
-- Company: USAFA/DFEC
-- Engineer: Silva
-- 
-- Create Date:    10:33:47 07/07/2012 
-- Design Name: 
-- Module Name:    MooreElevatorController_Silva - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: Code completed by C3C Demore, Mealy implementation of elevator FSM
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MealyElevatorController_Shell is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           stop : in  STD_LOGIC;
           up_down : in  STD_LOGIC;
           floor : out  STD_LOGIC_VECTOR (3 downto 0);
			  nextfloor : out std_logic_vector (3 downto 0));
end MealyElevatorController_Shell;

architecture Behavioral of MealyElevatorController_Shell is

type floor_state_type is (floor1, floor2, floor3, floor4);

signal current_state : floor_state_type;
signal next_state : floor_state_type;

begin

---------------------------------------------------------
--Code your Mealy machine next-state process below
--Question: Will it be different from your Moore Machine?
---------------------------------------------------------
next_state_process : process (current_state, up_down, stop)
begin
			case current_state is
				when floor1 =>
					if (up_down = '1' and stop = '0') then
						next_state <= floor2;
					else
						next_state <= floor1;
					end if;
				when floor2 =>
					if (up_down = '1' and stop = '0') then
						next_state <= floor3;
					elsif(up_down = '0' and stop = '0') then
						next_state <= floor1;
					else
						next_state <= floor2;
					end if;
				when floor3 =>
					if (up_down = '1' and stop = '0') then
						next_state <= floor4;
					elsif(up_down = '0' and stop = '0') then
						next_state <= floor2;
					else
						next_state <= floor3;
					end if;
				when floor4 =>
					if (up_down = '0' and stop = '0') then
						next_state <= floor3;
					else
						next_state <= floor4;
					end if;
				when others =>
					next_state <= floor1;
			end case;
end process;


-- state memory

	state_process : process (clk, reset) 
	begin						
		if (reset = '1') then
			current_state <= floor1;
		elsif (rising_edge (clk)) then
			current_state <= next_state;
		end if;
		
	end process;

-----------------------------------------------------------
--Code your Ouput Logic for your Mealy machine below
--Remember, now you have 2 outputs (floor and nextfloor)
-----------------------------------------------------------
floor <= "0001" when (current_state = floor1) else
			"0010" when (current_state = floor2) else
			"0011" when (current_state = floor3) else
			"0100" when (current_state = floor4) else
			"0001";

nextfloor <= 	"0001" when (next_state = floor1) else
					"0010" when (next_state = floor2) else
					"0011" when (next_state = floor3) else
					"0100" when (next_state = floor4) else
					"0001";

end Behavioral;

